LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY sub8 IS 
    PORT(
        A: IN UNSIGNED(7 DOWNTO 0);
        B: IN UNSIGNED(7 DOWNTO 0);
        C: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END sub8;

ARCHITECTURE dataflow OF sub8 IS
BEGIN
    C <= STD_LOGIC_VECTOR(("00000000" & A) - ("00000000" & B));
END dataflow;            